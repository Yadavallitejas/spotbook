** Profile: "SCHEMATIC1-hello4"  [ D:\ae lab\exp-1\rc shift-SCHEMATIC1-hello4.sim ] 

** Creating circuit file "rc shift-SCHEMATIC1-hello4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 20 100 1000mega
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rc shift-SCHEMATIC1.net" 


.END
